`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Universidad: TEC
// Ingenieros: Anthony Artavia - Diego Huertas - Justin Segura
// 
// Nombre del Módulo: binario_a_BCD
// Nombre del Proyecto: Algoritmo de Booth
// Descripción: Recibe el número binario resultante de la multiplicación y lo transforma a código BCD.
// 
//////////////////////////////////////////////////////////////////////////////////


module binario_a_BCD(

    );
endmodule
